library verilog;
use verilog.vl_types.all;
entity sim74138_vlg_vec_tst is
end sim74138_vlg_vec_tst;
