library verilog;
use verilog.vl_types.all;
entity chooser3_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end chooser3_vlg_check_tst;
