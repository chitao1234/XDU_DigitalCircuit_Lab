library verilog;
use verilog.vl_types.all;
entity async4_vlg_vec_tst is
end async4_vlg_vec_tst;
