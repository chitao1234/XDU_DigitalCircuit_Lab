library verilog;
use verilog.vl_types.all;
entity matrix_vlg_check_tst is
    port(
        COL1            : in     vl_logic;
        COL2            : in     vl_logic;
        COL3            : in     vl_logic;
        COL4            : in     vl_logic;
        COL5            : in     vl_logic;
        COL6            : in     vl_logic;
        COL7            : in     vl_logic;
        COL8            : in     vl_logic;
        ROW1            : in     vl_logic;
        ROW2            : in     vl_logic;
        ROW3            : in     vl_logic;
        ROW4            : in     vl_logic;
        ROW5            : in     vl_logic;
        ROW6            : in     vl_logic;
        ROW7            : in     vl_logic;
        ROW8            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end matrix_vlg_check_tst;
