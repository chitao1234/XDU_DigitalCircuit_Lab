library verilog;
use verilog.vl_types.all;
entity sim7483 is
    port(
        S1              : out    vl_logic;
        B4              : in     vl_logic;
        C0              : in     vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        A3              : in     vl_logic;
        B3              : in     vl_logic;
        A4              : in     vl_logic;
        S2              : out    vl_logic;
        S3              : out    vl_logic;
        S4              : out    vl_logic;
        C4              : out    vl_logic
    );
end sim7483;
