library verilog;
use verilog.vl_types.all;
entity sync4_vlg_vec_tst is
end sync4_vlg_vec_tst;
