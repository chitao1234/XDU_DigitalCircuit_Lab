library verilog;
use verilog.vl_types.all;
entity design4adder_vlg_vec_tst is
end design4adder_vlg_vec_tst;
