library verilog;
use verilog.vl_types.all;
entity mux41_vlg_vec_tst is
end mux41_vlg_vec_tst;
