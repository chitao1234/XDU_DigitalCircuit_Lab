library verilog;
use verilog.vl_types.all;
entity design24dec_vlg_sample_tst is
    port(
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        Ee              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end design24dec_vlg_sample_tst;
