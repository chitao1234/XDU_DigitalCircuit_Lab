library verilog;
use verilog.vl_types.all;
entity rssim_vlg_vec_tst is
end rssim_vlg_vec_tst;
