library verilog;
use verilog.vl_types.all;
entity chooser3_vlg_vec_tst is
end chooser3_vlg_vec_tst;
