library verilog;
use verilog.vl_types.all;
entity jksim_vlg_vec_tst is
end jksim_vlg_vec_tst;
