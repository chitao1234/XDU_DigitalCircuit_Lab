library verilog;
use verilog.vl_types.all;
entity sim7483_vlg_vec_tst is
end sim7483_vlg_vec_tst;
