library verilog;
use verilog.vl_types.all;
entity design24dec_vlg_vec_tst is
end design24dec_vlg_vec_tst;
